-- lcd1602.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lcd1602 is
	port (
		address     : in    std_logic                    := '0';             --   avalon_lcd_slave.address
		chipselect  : in    std_logic                    := '0';             --                   .chipselect
		read        : in    std_logic                    := '0';             --                   .read
		write       : in    std_logic                    := '0';             --                   .write
		writedata   : in    std_logic_vector(7 downto 0) := (others => '0'); --                   .writedata
		readdata    : out   std_logic_vector(7 downto 0);                    --                   .readdata
		waitrequest : out   std_logic;                                       --                   .waitrequest
		clk         : in    std_logic                    := '0';             --                clk.clk
		LCD_DATA    : inout std_logic_vector(7 downto 0) := (others => '0'); -- external_interface.DATA
		LCD_ON      : out   std_logic;                                       --                   .ON
		LCD_BLON    : out   std_logic;                                       --                   .BLON
		LCD_EN      : out   std_logic;                                       --                   .EN
		LCD_RS      : out   std_logic;                                       --                   .RS
		LCD_RW      : out   std_logic;                                       --                   .RW
		reset       : in    std_logic                    := '0'              --              reset.reset
	);
end entity lcd1602;

architecture rtl of lcd1602 is
	component lcd1602_character_lcd_0 is
		port (
			clk         : in    std_logic                    := 'X';             -- clk
			reset       : in    std_logic                    := 'X';             -- reset
			address     : in    std_logic                    := 'X';             -- address
			chipselect  : in    std_logic                    := 'X';             -- chipselect
			read        : in    std_logic                    := 'X';             -- read
			write       : in    std_logic                    := 'X';             -- write
			writedata   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(7 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                       -- waitrequest
			LCD_DATA    : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_ON      : out   std_logic;                                       -- export
			LCD_BLON    : out   std_logic;                                       -- export
			LCD_EN      : out   std_logic;                                       -- export
			LCD_RS      : out   std_logic;                                       -- export
			LCD_RW      : out   std_logic                                        -- export
		);
	end component lcd1602_character_lcd_0;

begin

	character_lcd_0 : component lcd1602_character_lcd_0
		port map (
			clk         => clk,         --                clk.clk
			reset       => reset,       --              reset.reset
			address     => address,     --   avalon_lcd_slave.address
			chipselect  => chipselect,  --                   .chipselect
			read        => read,        --                   .read
			write       => write,       --                   .write
			writedata   => writedata,   --                   .writedata
			readdata    => readdata,    --                   .readdata
			waitrequest => waitrequest, --                   .waitrequest
			LCD_DATA    => LCD_DATA,    -- external_interface.export
			LCD_ON      => LCD_ON,      --                   .export
			LCD_BLON    => LCD_BLON,    --                   .export
			LCD_EN      => LCD_EN,      --                   .export
			LCD_RS      => LCD_RS,      --                   .export
			LCD_RW      => LCD_RW       --                   .export
		);

end architecture rtl; -- of lcd1602
